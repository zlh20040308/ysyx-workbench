module ysyx_23060337_EXU(
    input clk,
    input [31:0] rd,
    input [31:0] rs1,
    input [31:0] rs2,
    input [31:0] imm,
    input [2:0] funct3,
    input [6:0] funct7,
    input [6:0] opcode
);




endmodule