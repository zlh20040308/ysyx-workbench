module example();
endmodule
