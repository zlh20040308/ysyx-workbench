module ysyx_23060337_EXU(
    input clk,
    input rst,
    input [31:0] inst,
    output reg [31:0] pc,
);




endmodule