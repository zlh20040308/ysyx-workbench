module ysyx_23060337_IFU(
    input clk,
    input rst,
    input reg [31:0] pc,
    output reg [31:0] inst,
);




endmodule